VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ws_ip__credits
  CLASS BLOCK ;
  FOREIGN gf180mcu_ws_ip__credits ;
  ORIGIN 0.000 0.000 ;
  SIZE 143.25 BY 143.25 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 143.25 143.25 ;
  END
END gf180mcu_ws_ip__credits
END LIBRARY

