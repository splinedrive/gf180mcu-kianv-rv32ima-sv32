module gf180mcu_ws_ip__credits;
endmodule
